library verilog;
use verilog.vl_types.all;
entity maxpool_tb is
end maxpool_tb;
