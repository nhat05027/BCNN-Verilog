library verilog;
use verilog.vl_types.all;
entity tb_FullyConnect is
end tb_FullyConnect;
