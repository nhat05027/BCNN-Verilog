library verilog;
use verilog.vl_types.all;
entity tb_conv is
end tb_conv;
