library verilog;
use verilog.vl_types.all;
entity bnorm_tb is
end bnorm_tb;
