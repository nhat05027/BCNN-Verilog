//Copyright (C)2014-2024 Gowin Semiconductor Corporation.
//All rights reserved.
//File Title: IP file
//Tool Version: V1.9.10.03 Education (64-bit)
//Part Number: GW1NR-LV9QN88PC6/I5
//Device: GW1NR-9
//Device Version: C
//Created Time: Thu Apr 17 17:19:05 2025

module Gowin_SDPB (dout, clka, cea, reseta, clkb, ceb, resetb, oce, ada, din, adb);

output [7:0] dout;
input clka;
input cea;
input reseta;
input clkb;
input ceb;
input resetb;
input oce;
input [9:0] ada;
input [7:0] din;
input [9:0] adb;

wire [23:0] sdpb_inst_0_dout_w;
wire gw_gnd;

assign gw_gnd = 1'b0;

SDPB sdpb_inst_0 (
    .DO({sdpb_inst_0_dout_w[23:0],dout[7:0]}),
    .CLKA(clka),
    .CEA(cea),
    .RESETA(reseta),
    .CLKB(clkb),
    .CEB(ceb),
    .RESETB(resetb),
    .OCE(oce),
    .BLKSELA({gw_gnd,gw_gnd,gw_gnd}),
    .BLKSELB({gw_gnd,gw_gnd,gw_gnd}),
    .ADA({gw_gnd,ada[9:0],gw_gnd,gw_gnd,gw_gnd}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[7:0]}),
    .ADB({gw_gnd,adb[9:0],gw_gnd,gw_gnd,gw_gnd})
);

defparam sdpb_inst_0.READ_MODE = 1'b0;
defparam sdpb_inst_0.BIT_WIDTH_0 = 8;
defparam sdpb_inst_0.BIT_WIDTH_1 = 8;
defparam sdpb_inst_0.BLK_SEL_0 = 3'b000;
defparam sdpb_inst_0.BLK_SEL_1 = 3'b000;
defparam sdpb_inst_0.RESET_MODE = "SYNC";
defparam sdpb_inst_0.INIT_RAM_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_0.INIT_RAM_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_0.INIT_RAM_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_0.INIT_RAM_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_0.INIT_RAM_04 = 256'h4600000000000000E03200000000000000000000000000000000000000000000;
defparam sdpb_inst_0.INIT_RAM_05 = 256'h000000A89400000000000000E77900000000000000000000000000000000001D;
defparam sdpb_inst_0.INIT_RAM_06 = 256'h0000000000000BD26000000000000000E7C30400000000000000000000000000;
defparam sdpb_inst_0.INIT_RAM_07 = 256'h0000000000000000000015FC720000000000000086FC45000000000000000000;
defparam sdpb_inst_0.INIT_RAM_08 = 256'h000000000000000000000000000015FCC0000000000000000CD9EC2D00000000;
defparam sdpb_inst_0.INIT_RAM_09 = 256'h0000D3F2540000000000000000000000000015FDFF120000000000000035F7A8;
defparam sdpb_inst_0.INIT_RAM_0A = 256'h0000000000006AFCA90000000000000000000000000005BDFD8D000000000000;
defparam sdpb_inst_0.INIT_RAM_0B = 256'hD3FC860000000000000000FCE10F0000000000000000000000000042FAE82000;
defparam sdpb_inst_0.INIT_RAM_0C = 256'h00000000A7FCA90000000000000000A4FC160000000000000000000000000000;
defparam sdpb_inst_0.INIT_RAM_0D = 256'h00000000000000006BFDFD1600000000000012D1CC0900000000000000000000;
defparam sdpb_inst_0.INIT_RAM_0E = 256'h0000000000000000000000006AFCFCC3A48155555555C7FCA900000000000000;
defparam sdpb_inst_0.INIT_RAM_0F = 256'h0000000000000000000000000000000009FCFCFBE7E8FCFCFCFCF5AA29000000;
defparam sdpb_inst_0.INIT_RAM_10 = 256'h000000000000000000000000000000000000000000FCFCA10000545454543100;
defparam sdpb_inst_0.INIT_RAM_11 = 256'h0000000000000000000000000000000000000000000000002DFCFC7F00000000;
defparam sdpb_inst_0.INIT_RAM_12 = 256'h00FCFC7F00000000000000000000000000000000000000000000000000FDFD80;
defparam sdpb_inst_0.INIT_RAM_13 = 256'h0000000000F4FC87000000000000000000000000000000000000000000000000;
defparam sdpb_inst_0.INIT_RAM_14 = 256'h0000000000000000006FECE80000000000000000000000000000000000000000;
defparam sdpb_inst_0.INIT_RAM_15 = 256'h000000000000000000000000000042B300000000000000000000000000000000;
defparam sdpb_inst_0.INIT_RAM_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_0.INIT_RAM_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sdpb_inst_0.INIT_RAM_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;

endmodule //Gowin_SDPB
