library verilog;
use verilog.vl_types.all;
entity tb_cnn_data is
end tb_cnn_data;
