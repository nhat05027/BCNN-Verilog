library verilog;
use verilog.vl_types.all;
entity tb_cnn is
end tb_cnn;
